-- router module
-- forwards packets to neighbouring routers and local network adapter
-- routing priorities given to : local, N, E, S, W inputs
-- each input has 2 levels of buffers
-- packets held in buffers when a higher priority input also wants to write to same output
-- also held in buffers if the output is busy
-- an output is set to busy when the input buffer is being used and therefore cannot take any more input packets

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity router is
	generic (
		node_ID 	: std_logic_vector(3 downto 0)
	);
	port (
		clk     	: in std_logic;
		nreset	: in std_logic;
		
		--busy signals 		- 0 = local, 1 = north, 2 = east, 3 = south, 4 = west
		busy_in 			: in std_logic_vector(4 downto 0);
		busy_out 		: out std_logic_vector(4 downto 0);

		local_pkt_in 	: in std_logic_vector(48 downto 0);
		local_pkt_out 	: out std_logic_vector(48 downto 0);
		
		north_pkt_in 	: in std_logic_vector(48 downto 0);
		north_pkt_out 	: out std_logic_vector(48 downto 0);
		
		east_pkt_in 	: in std_logic_vector(48 downto 0);
		east_pkt_out 	: out std_logic_vector(48 downto 0);
		
		south_pkt_in 	: in std_logic_vector(48 downto 0);
		south_pkt_out 	: out std_logic_vector(48 downto 0);
		
		west_pkt_in 	: in std_logic_vector(48 downto 0);
		west_pkt_out 	: out std_logic_vector(48 downto 0)
		
	);
end router;

architecture rtl of router is

	-- bus_array - 0 = local, 1 = north, 2 = east, 3 = south, 4 = west
	type bus_array_type is array(integer range 4 downto 0) of std_logic_vector(48 downto 0);

--	signal bus_array_in 			: bus_array_type;
	signal bus_array_boundary_in 		: bus_array_type;
	signal bus_array_out 			: bus_array_type;



	signal buffer_level1 			: bus_array_type;
	signal buffer_level2 			: bus_array_type;
		
	signal buffer_level1_used 		: std_logic_vector(4 downto 0) := "00000";
	signal buffer_level2_used 		: std_logic_vector(4 downto 0) := "00000";
	
begin

	bus_array_boundary_in(0) <= local_pkt_in;
	bus_array_boundary_in(1) <= north_pkt_in;
	bus_array_boundary_in(2) <= east_pkt_in;
	bus_array_boundary_in(3) <= south_pkt_in;
	bus_array_boundary_in(4) <= west_pkt_in;
		
	local_pkt_out 	<= bus_array_out(0);
	north_pkt_out 	<= bus_array_out(1);
	east_pkt_out 	<= bus_array_out(2);
	south_pkt_out 	<= bus_array_out(3);
	west_pkt_out 	<= bus_array_out(4);
	
	busy_out		<= buffer_level1_used;
		
	process(clk)
		variable is_collision 	: std_logic_vector(4 downto 0); 
		
		type bus_array_type is array(integer range 4 downto 0) of std_logic_vector(48 downto 0);
		
		variable bus_array_in 			: bus_array_type;
		
		type yx_array_type is array(integer range 4 downto 0) of std_logic_vector(1 downto 0);
		
		variable y 					: yx_array_type;	
		variable x 					: yx_array_type;
	
		variable sign_y 				: std_logic_vector(4 downto 0);	
		variable sign_x 				: std_logic_vector(4 downto 0);

		type integer_array_type is array(integer range 4 downto 0) of natural range 0 to 6;
		variable direction 			: integer_array_type;
		
	begin
			
		if (rising_edge(clk)) then 
			if nreset = '0' then
				bus_array_out(0) <= (others => '0');
				bus_array_out(1) <= (others => '0');
				bus_array_out(2) <= (others => '0');
				bus_array_out(3) <= (others => '0');
				bus_array_out(4) <= (others => '0');
				
				buffer_level1_used <= "00000";
				buffer_level2_used <= "00000";
				
				buffer_level1(0) <= (others => '0');
				buffer_level1(1) <= (others => '0');
				buffer_level1(2) <= (others => '0');
				buffer_level1(3) <= (others => '0');
				buffer_level1(4) <= (others => '0');
				
				buffer_level2(0) <= (others => '0');
				buffer_level2(1) <= (others => '0');
				buffer_level2(2) <= (others => '0');
				buffer_level2(3) <= (others => '0');
				buffer_level2(4) <= (others => '0');
				
			else
				--default values
				bus_array_out(0) <= (others => '0');
				bus_array_out(1) <= (others => '0');
				bus_array_out(2) <= (others => '0');
				bus_array_out(3) <= (others => '0');
				bus_array_out(4) <= (others => '0');

			
				for i in 0 to 4 loop --for each input bus array
					
					-- choose an input (packet_in or buffer1)
					if (buffer_level1_used(i) = '1' ) then
						bus_array_in(i) := buffer_level1(i);
					else
						bus_array_in(i) := bus_array_boundary_in(i);
					end if;
					
					sign_y(i) := bus_array_in(i)(48);
					sign_x(i) := bus_array_in(i)(45);
					y(i) := bus_array_in(i)(47 downto 46);
					x(i) := bus_array_in(i)(44 downto 43);
					
					--calculate desired direction
					if ((bus_array_in(i)(42) = '0' and bus_array_in(i)(41) = '0' and bus_array_in(i)(40) = '0')) then
						direction(i) := 6; --empty
					elsif (y(i) /= "00") then
						if (sign_y(i) = '1') then
							direction(i) := 1; --north
						elsif (sign_y(i) = '0') then
							direction(i) := 3; --south
						end if;
					elsif (x(i) /= "00") then
						if (sign_x(i) = '1') then
							direction(i) := 4; --west
						elsif (sign_x(i) = '0') then
							direction(i) := 2; --east
						end if;
					elsif (y(i) = "00" and x(i) = "00") then
						direction(i) := 0; --local
					end if;				
					
					--if not empty packet
					if(bus_array_in(i)(42) = '1' or bus_array_in(i)(41) = '1' or bus_array_in(i)(40) = '1') then

						--check for collisions with busy_in and all previous bus_array_in's

						is_collision(i) := '0'; --flag

						if( busy_in(direction(i)) = '1') then --check busy signal
							is_collision(i) := '1';
						elsif( i > 0 ) then
							--check bus_array_in's with higher priority
							for j in 0 to i-1 loop 
								if(direction(i) = direction(j)) then --this does not include if they're both empty due to outer if statement above
									is_collision(i) := '1';
								end if;
							end loop;

						end if;
					
						if (buffer_level1_used(i) = '1' and is_collision(i) = '1') then
							buffer_level1(i) <= buffer_level1(i);
							buffer_level1_used(i) <= '1';
						elsif (buffer_level1_used(i) = '1' and buffer_level2_used(i) ='1' and is_collision(i) = '0') then
							buffer_level1(i) <= buffer_level2(i);
							buffer_level1_used(i) <= '1';
						elsif ((bus_array_boundary_in(i)(42) = '1' or bus_array_boundary_in(i)(41) = '1' or bus_array_boundary_in(i)(40) = '1')
									and buffer_level1_used(i) = '1' and buffer_level2_used(i) ='0' and is_collision(i) = '0') then
							
							buffer_level1(i) <= bus_array_boundary_in(i);
							buffer_level1_used(i) <= '1';
						elsif ((bus_array_boundary_in(i)(42) = '1' or bus_array_boundary_in(i)(41) = '1' or bus_array_boundary_in(i)(40) = '1')
									and buffer_level1_used(i) = '0' and buffer_level2_used(i) ='0' and is_collision(i) = '1') then
							
							buffer_level1(i) <= bus_array_boundary_in(i);
							buffer_level1_used(i) <= '1';
						else
							buffer_level1(i) <= (others => '0');
							buffer_level1_used(i) <= '0';
						end if;
						
						if (buffer_level1_used(i) = '1' and buffer_level2_used(i) = '1' and is_collision(i) = '1') then
							buffer_level2(i) <= buffer_level2(i);
							buffer_level2_used(i) <= '1';
						elsif ((bus_array_boundary_in(i)(42) = '1' or bus_array_boundary_in(i)(41) = '1' or bus_array_boundary_in(i)(40) = '1') 
								and buffer_level1_used(i) = '1' and buffer_level2_used(i) = '1' and is_collision(i) = '0') then
							
							buffer_level2(i) <= bus_array_boundary_in(i);
							buffer_level2_used(i) <= '1';
						elsif ((bus_array_boundary_in(i)(42) = '1' or bus_array_boundary_in(i)(41) = '1' or bus_array_boundary_in(i)(40) = '1') 
								and buffer_level1_used(i) = '1' and buffer_level2_used(i) = '0' and is_collision(i) = '1') then
								
							buffer_level2(i) <= bus_array_boundary_in(i);
							buffer_level2_used(i) <= '1';
						else
							buffer_level2(i) <= (others => '0');
							buffer_level2_used(i) <= '0';
						end if;			
							

						--send to output
						if (is_collision(i) = '0') then
							
							if (y(i) /= "00") then
								if (sign_y(i) = '1') then
									bus_array_out(1) <= sign_y(i) & std_logic_vector(unsigned(y(i)) - 1) & sign_x(i) & x(i) & bus_array_in(i)(42 downto 0);
								elsif (sign_y(i) = '0') then
									bus_array_out(3) <= sign_y(i) & std_logic_vector(unsigned(y(i)) - 1) & sign_x(i) & x(i) & bus_array_in(i)(42 downto 0);
								end if;
							elsif (x(i) /= "00") then
								if (sign_x(i) = '1') then
									bus_array_out(4) <= sign_y(i) & y(i) & sign_x(i) & std_logic_vector(unsigned(x(i)) - 1) & bus_array_in(i)(42 downto 0);
								elsif (sign_x(i) = '0') then
									bus_array_out(2) <= sign_y(i) & y(i) & sign_x(i) & std_logic_vector(unsigned(x(i)) - 1) & bus_array_in(i)(42 downto 0);
								end if;
							elsif (y(i) = "00" and x(i) = "00") then
								bus_array_out(0) <= bus_array_in(i); -- destination node reached, to local
							end if;
						
						end if; --is collision
					end if; 	--empty packet
				end loop;		--i	
			end if; 			--reset
		end if; 				--rising_edge clk
				
	end process;

end rtl;

